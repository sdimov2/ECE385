module note_rom ( input [5:0]	addr,
						output [48:0]	data
					 );

	parameter ADDR_WIDTH = 6;
   parameter DATA_WIDTH =  49;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {

			49'h000001FF00000, // 0
			49'h000001FF00000,
			49'h000001FF00000,
			49'h000001FF00000,
			49'h0000000000000,
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,
			49'h0000000000000,
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,
			49'h0000000000000,
			49'h0000000000000,
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,
			49'h0000000000000,
			49'h0000000000000,
			49'h0000000000000,
			49'h0000000000000,
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,			
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,
			49'h0000000000000,
			49'h0000000000000,
			49'h0000000000000,
			49'h0000000000000,
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,
			49'h0000000000000,
			49'h0000000000000,
			49'hFFFFFFFFFFFFF,
			49'hFFFFFFFFFFFFF,
			49'h0000000000000,
			49'h000001FF00000,
			49'h000001FF00000,
			49'h000001FF00000,
			49'h000001FF00000

        };

	assign data = ROM[addr];

endmodule  