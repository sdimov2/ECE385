module I2S_interface 
(
	input 	I2S_DIN,
	output 	I2S_DOUT,
	output	LRCLK,
	output	SCLK
);


endmodule