module fpga_guitar_hero(

      ///////// Clocks /////////
      input    MAX10_CLK1_50,

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,





      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N,
		input					 A2,
		input					 A3,
		input					 A4
);

logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST;
logic I2C_SCL_IN, I2C_SCL_OUT, I2C_SDA_IN, I2C_SDA_OUT;
logic I2S_LRCLK, I2S_MCLK, I2S_DOUT, I2S_DIN;
logic [3:0] hex_num_4, hex_num_3, hex_num_1, hex_num_0; //4 bit input hex digits
logic [1:0] signs;
logic [1:0] hundreds;

assign ARDUINO_IO[10] = SPI0_CS_N;
assign ARDUINO_IO[13] = SPI0_SCLK;
assign ARDUINO_IO[11] = SPI0_MOSI;
assign ARDUINO_IO[12] = 1'bZ;
assign SPI0_MISO = ARDUINO_IO[12];

assign ARDUINO_IO[3] = I2S_MCLK;
assign ARDUINO_IO[1] = I2S_DOUT;

assign ARDUINO_IO[14] = I2C_SDA_OUT ? 1'b0 : 1'bz;
assign ARDUINO_IO[15] = I2C_SCL_OUT ? 1'b0 : 1'bz;

assign I2C_SDA_IN = ARDUINO_IO[14];
assign I2C_SCL_IN = ARDUINO_IO[15];

//Assignments specific to Circuits At Home UHS_20
assign ARDUINO_RESET_N = USB_RST;
assign ARDUINO_IO[7] = USB_RST;//USB reset 
assign ARDUINO_IO[8] = 1'bZ; //this is GPX (set to input)
assign USB_GPX = 1'b0;//GPX is not needed for standard USB host - set to 0 to prevent interrupt


//Assign uSD CS to '1' to prevent uSD card from interfering with USB Host (if uSD card is plugged in)
assign ARDUINO_IO[6] = 1'b1;

//HEX drivers to convert numbers to HEX output
HexDriver hex_driver4 (hex_num_4, HEX4[6:0]);
assign HEX4[7] = 1'b1;

HexDriver hex_driver3 (hex_num_3, HEX3[6:0]);
assign HEX3[7] = 1'b1;

HexDriver hex_driver1 (hex_num_1, HEX1[6:0]);
assign HEX1[7] = 1'b1;

HexDriver hex_driver0 (hex_num_0, HEX0[6:0]);
assign HEX0[7] = 1'b1;

//fill in the hundreds digit as well as the negative sign
assign HEX5 = {1'b1, ~signs[1], 3'b111, ~hundreds[1], ~hundreds[1], 1'b1};
assign HEX2 = {1'b1, ~signs[0], 3'b111, ~hundreds[0], ~hundreds[0], 1'b1};
	
logic [1:0] clkdiv;

always @(posedge MAX10_CLK1_50) begin
	if (clkdiv == 2'b0)
		I2S_MCLK <= ~I2S_MCLK;
	clkdiv <= clkdiv + 1;
end

fpga_guitar_hero_soc u0 (
		.clk_clk                           (MAX10_CLK1_50),    //clk.clk
		.reset_reset_n                     (1'b1),             //reset.reset_n

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),            				   //clk_sdram.clk
	   .sdram_wire_addr(DRAM_ADDR),               			   //sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),                			   //.ba
		.sdram_wire_cas_n(DRAM_CAS_N),              		   //.cas_n
		.sdram_wire_cke(DRAM_CKE),                 			   //.cke
		.sdram_wire_cs_n(DRAM_CS_N),                		   //.cs_n
		.sdram_wire_dq(DRAM_DQ),                  			   //.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),                //.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),              		   //.ras_n
		.sdram_wire_we_n(DRAM_WE_N),                		   //.we_n
		

		.vga_red(VGA_R),          //        vga.red
		.vga_green(VGA_G),        //           .green
		.vga_blue(VGA_B),         //           .blue
		.vga_hs(VGA_HS),           //           .hs
		.vga_vs(VGA_VS),            //           .vs
		
		.spi_0_external_MISO(SPI0_MISO),     //   spi_0_external.MISO
		.spi_0_external_MOSI(SPI0_MOSI),     //                 .MOSI
		.spi_0_external_SCLK(SPI0_SCLK),     //                 .SCLK
		.spi_0_external_SS_n(SPI0_CSP_N),     //                 .SS_n
		
		.usb_gpx_export(USB_GPX),          //          usb_gpx.export
		.usb_irq_export(USB_IRQ),          //          usb_irq.export
		.usb_rst_export(USB_RST),          //          usb_rst.export
		
		.i2c_0_i2c_serial_sda_in(I2C_SDA_IN), // i2c_0_i2c_serial.sda_in
		.i2c_0_i2c_serial_scl_in(I2C_SCL_IN), //                 .scl_in
		.i2c_0_i2c_serial_sda_oe(I2C_SDA_OUT), //                 .sda_oe
		.i2c_0_i2c_serial_scl_oe(I2C_SCL_OUT), //                 .scl_oe
		
		.hex_digits_wire_export({hex_num_4, hex_num_3, hex_num_1, hex_num_0}),  //  hex_digits_wire.export
		.leds_wire_export({hundreds, signs, LEDR}),        //        leds_wire.export
		.frets_pio_wire_export({~A4, ~KEY[0], ~KEY[1], ~A3, ~A2})
	 );

endmodule
